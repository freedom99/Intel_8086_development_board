-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Thursday, October 16, 2014 20:33:36 Bangladesh Standard Time

